[[.tagcollection ]]

[[.begin name=boxlet singleton=True ]]
[[.attr name=width default=300 ]]
[[.attr name=lines default=5 ]]

[[.import names="pool"]] [[-- creates pool alias for serverglobals --]]

[[--
  You can and often should put the handlers in a separate file,
  with the class it associates with where applicable.  Here
  We just inline our handler; for an example of the other,
  see the to-do demo.
--]]
[[!
def chatbox_addline(self, api, newline):
    # (use setdefault() in case server restarted)
    api.pool.setdefault('chatlines', []).append(newline)
    api.pool['chatlines'] = api.pool['chatlines'][:100] # remembers max of 100
]]

<div width="[[= width ]]">
  [[\
     i = -int(lines)
     line = None # for first export
  ]]
  [[ for line in pool.setdefault('chatlines', [])[i:]:{ ]]
  <div>[[= line ]]</div>
  [[ } ]]
  <div>
  <f:text name=newline value="" />
  <f:submit handler='self.chatbox_addline' value="Send" />
  <f:submit value="Refresh" />
  </div>
</div>

[[.export var=line as=last ]] [[-- sends this variable to the calling scope --]]
[[.end]]
