[[.begin name=bold buffers=True]]

<b>[[=_contents]]</b>

[[.end]]